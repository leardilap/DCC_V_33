LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DCC_V_33_TB IS
END DCC_V_33_TB;

ARCHITECTURE DCC_V_33_TB_ARCH OF DCC_V_33_TB IS

    COMPONENT DCC_V_33 IS
        PORT (
			OSC_50 			: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			
			--//////// LED //////////
			LEDG			: OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
			LEDR			: OUT STD_LOGIC_VECTOR (17 DOWNTO 0);

			--//////// KEY //////////
			KEY				: IN STD_LOGIC_VECTOR (3 DOWNTO 0);

			--//////// SW //////////
			SW				: IN STD_LOGIC_VECTOR (17 DOWNTO 0);

			--//////// HSMC //////////
			AD_SCLK			: IN STD_LOGIC;
			AD_SDIO			: IN STD_LOGIC;
			ADA_D			: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
			ADA_DCO			: IN STD_LOGIC;
			ADA_OE			: OUT STD_LOGIC;
			ADA_OR			: IN STD_LOGIC;
			ADA_SPI_CS		: OUT STD_LOGIC;
			ADB_D			: IN STD_LOGIC_VECTOR (13 DOWNTO 0);
			ADB_DCO			: IN STD_LOGIC;
			ADB_OE			: OUT STD_LOGIC;
			ADB_OR			: IN STD_LOGIC;
			ADB_SPI_CS		: OUT STD_LOGIC;
			AIC_BCLK		: IN STD_LOGIC;
			AIC_DIN			: OUT STD_LOGIC;
			AIC_DOUT		: IN STD_LOGIC;
			AIC_LRCIN		: IN STD_LOGIC;
			AIC_LRCOUT		: IN STD_LOGIC;
			AIC_SPI_CS		: OUT STD_LOGIC;
			AIC_XCLK		: OUT STD_LOGIC;
			CLKIN1			: IN STD_LOGIC;
			CLKOUT0			: OUT STD_LOGIC;
			DA				: OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
			DB				: OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
			FPGA_CLK_A_N	: OUT STD_LOGIC;
			FPGA_CLK_A_P	: OUT STD_LOGIC;
			FPGA_CLK_B_N	: OUT STD_LOGIC;
			FPGA_CLK_B_P	: OUT STD_LOGIC;
			J1_152			: IN STD_LOGIC;
			XT_IN_N			: IN STD_LOGIC;
			XT_IN_P 		: IN STD_LOGIC
		);
    END COMPONENT DCC_V_33;

	SIGNAL		OSC_50 			: STD_LOGIC_VECTOR (2 DOWNTO 0);
			
	--//////// LED //////
	SIGNAL		LEDG			: STD_LOGIC_VECTOR (8 DOWNTO 0);
	SIGNAL		LEDR			: STD_LOGIC_VECTOR (17 DOWNTO 0);
    
	--//////// KEY //////
	SIGNAL		KEY				: STD_LOGIC_VECTOR (3 DOWNTO 0);
    
	--//////// SW //////
	SIGNAL		SW				: STD_LOGIC_VECTOR (17 DOWNTO 0);
    
	--//////// HSMC //////
	SIGNAL		AD_SCLK			: STD_LOGIC;
	SIGNAL		AD_SDIO			: STD_LOGIC;
	SIGNAL		ADA_D			: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL		ADA_DCO			: STD_LOGIC;
	SIGNAL		ADA_OE			: STD_LOGIC;
	SIGNAL		ADA_OR			: STD_LOGIC;
	SIGNAL		ADA_SPI_CS		: STD_LOGIC;
	SIGNAL		ADB_D			: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL		ADB_DCO			: STD_LOGIC;
	SIGNAL		ADB_OE			: STD_LOGIC;
	SIGNAL		ADB_OR			: STD_LOGIC;
	SIGNAL		ADB_SPI_CS		: STD_LOGIC;
	SIGNAL		AIC_BCLK		: STD_LOGIC;
	SIGNAL		AIC_DIN			: STD_LOGIC;
	SIGNAL		AIC_DOUT		: STD_LOGIC;
	SIGNAL		AIC_LRCIN		: STD_LOGIC;
	SIGNAL		AIC_LRCOUT		: STD_LOGIC;
	SIGNAL		AIC_SPI_CS		: STD_LOGIC;
	SIGNAL		AIC_XCLK		: STD_LOGIC;
	SIGNAL		CLKIN1			: STD_LOGIC;
	SIGNAL		CLKOUT0			: STD_LOGIC;
	SIGNAL		DA				: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL		DB				: STD_LOGIC_VECTOR (13 DOWNTO 0);
	SIGNAL		FPGA_CLK_A_N	: STD_LOGIC;
	SIGNAL		FPGA_CLK_A_P	: STD_LOGIC;
	SIGNAL		FPGA_CLK_B_N	: STD_LOGIC;
	SIGNAL		FPGA_CLK_B_P	: STD_LOGIC;
	SIGNAL		J1_152			: STD_LOGIC;
	SIGNAL		XT_IN_N			: STD_LOGIC;
	SIGNAL		XT_IN_P 		: STD_LOGIC;

    CONSTANT OSC_50_Period : TIME := 20 ns;
	
BEGIN
	
	UUT_DCC_V_33 : DCC_V_33
        PORT MAP(
			OSC_50 			  => OSC_50,
			LEDG			  => LEDG,			
			LEDR			  => LEDR,			
			KEY				  => KEY,			
			SW				  => SW,	
			AD_SCLK			  => AD_SCLK,			
			AD_SDIO			  => AD_SDIO,			
			ADA_D			  => ADA_D,			
			ADA_DCO			  => ADA_DCO,			
			ADA_OE			  => ADA_OE,			
			ADA_OR			  => ADA_OR,			
			ADA_SPI_CS		  => ADA_SPI_CS,		
			ADB_D			  => ADB_D,			
			ADB_DCO			  => ADB_DCO,			
			ADB_OE			  => ADB_OE,			
			ADB_OR			  => ADB_OR,			
			ADB_SPI_CS		  => ADB_SPI_CS,	
			AIC_BCLK		  => AIC_BCLK,		
			AIC_DIN			  => AIC_DIN,			
			AIC_DOUT		  => AIC_DOUT,		
			AIC_LRCIN		  => AIC_LRCIN,		
			AIC_LRCOUT		  => AIC_LRCOUT,		
			AIC_SPI_CS		  => AIC_SPI_CS,		
			AIC_XCLK		  => AIC_XCLK,		
			CLKIN1			  => CLKIN1,			
			CLKOUT0			  => CLKOUT0,			
			DA				  => DA,				
			DB				  => DB,				
			FPGA_CLK_A_N	  => FPGA_CLK_A_N,	
			FPGA_CLK_A_P	  => FPGA_CLK_A_P,	
			FPGA_CLK_B_N	  => FPGA_CLK_B_N,	
			FPGA_CLK_B_P	  => FPGA_CLK_B_P,	
			J1_152			  => J1_152,			
			XT_IN_N			  => XT_IN_N,			
			XT_IN_P 		  => XT_IN_P 		
		);
	
	OSC_50(0) <= NOT OSC_50(0) AFTER OSC_50_Period/2;
	KEY(3) <= '1';
	ADA_DCO <= OSC_50(0);
	ADB_DCO <= OSC_50(0);
	
	ADB_D	<= STD_LOGIC_VECTOR( TO_UNSIGNED(215, 14) );
	ADB_D	<= STD_LOGIC_VECTOR( TO_UNSIGNED(1215, 14) );
	
END DCC_V_33_TB_ARCH;